library verilog;
use verilog.vl_types.all;
entity menor_vlg_vec_tst is
end menor_vlg_vec_tst;
