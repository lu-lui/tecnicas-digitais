library verilog;
use verilog.vl_types.all;
entity tdexemplo5_vlg_vec_tst is
end tdexemplo5_vlg_vec_tst;
