library verilog;
use verilog.vl_types.all;
entity display_mux_vlg_vec_tst is
end display_mux_vlg_vec_tst;
