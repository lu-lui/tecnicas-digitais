library verilog;
use verilog.vl_types.all;
entity subtrator4bits_vlg_vec_tst is
end subtrator4bits_vlg_vec_tst;
