library verilog;
use verilog.vl_types.all;
entity sr_b_vlg_vec_tst is
end sr_b_vlg_vec_tst;
