library verilog;
use verilog.vl_types.all;
entity tdexemplo5 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        S               : out    vl_logic
    );
end tdexemplo5;
