library verilog;
use verilog.vl_types.all;
entity meio_somador_vlg_vec_tst is
end meio_somador_vlg_vec_tst;
