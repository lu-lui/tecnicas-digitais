library verilog;
use verilog.vl_types.all;
entity cod_bin_hexa_vlg_vec_tst is
end cod_bin_hexa_vlg_vec_tst;
