library verilog;
use verilog.vl_types.all;
entity multiplicador4bits_vlg_vec_tst is
end multiplicador4bits_vlg_vec_tst;
