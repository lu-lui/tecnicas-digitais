LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY seg7_somador IS
	PORT( 
		a, b :in std_logic_vector (3 downto 0);
		s: out std_logic_vector(6 downto 0);
		c4: out std_logic
		);
end seg7_somador;
architecture arq_seg7_somador of seg7_somador is
	SIGNAL n: std_logic_vector(3 downto 0);
	
	COMPONENT somador4bits
		PORT( 
		a, b :in std_logic_vector (3 downto 0);
		s:out std_logic_vector(3 downto 0);
		c4: out std_logic
		);
	END COMPONENT;
	
	COMPONENT seg7
		PORT( 
		entrada :in std_logic_vector(3 downto 0);
		s :out std_logic_vector (6 downto 0)
		);
	END COMPONENT;
	
	begin 
		somador: somador4bits
			port map (a => a, b => b, s => n, c4 => c4);
			
		segmento7: seg7
			port map (entrada => n, s => s);
			
	end arq_seg7_somador;
	