library verilog;
use verilog.vl_types.all;
entity tdexemplo5_vlg_check_tst is
    port(
        S               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end tdexemplo5_vlg_check_tst;
