library verilog;
use verilog.vl_types.all;
entity tdexemplo9_vlg_vec_tst is
end tdexemplo9_vlg_vec_tst;
