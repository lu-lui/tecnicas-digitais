library verilog;
use verilog.vl_types.all;
entity somador4bits_vlg_vec_tst is
end somador4bits_vlg_vec_tst;
