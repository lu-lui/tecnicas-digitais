library verilog;
use verilog.vl_types.all;
entity a_xor_b_vlg_vec_tst is
end a_xor_b_vlg_vec_tst;
