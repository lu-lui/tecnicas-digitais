library verilog;
use verilog.vl_types.all;
entity sl_a_vlg_vec_tst is
end sl_a_vlg_vec_tst;
