library verilog;
use verilog.vl_types.all;
entity display_7seg_vlg_vec_tst is
end display_7seg_vlg_vec_tst;
