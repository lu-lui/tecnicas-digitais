library verilog;
use verilog.vl_types.all;
entity display_mult_vlg_vec_tst is
end display_mult_vlg_vec_tst;
