library verilog;
use verilog.vl_types.all;
entity meio_somador_vlg_check_tst is
    port(
        c_out           : in     vl_logic;
        s               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end meio_somador_vlg_check_tst;
